/////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//  NAME      :- Pradip Prajapati
//  FILE_NAME :- ahb_defines.svh
//  EDITED_BY :- Rajvi Padaria
//
//////////////////////////////////////////////////////////////////////////////////////////////////////////

`define ADDR_WIDTH 32
`define DATA_WIDTH 1024

