typedef uvm_sequencer#(apb_uart_tx)apb_uart_sqr; 
