//////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//  NAME      :- Pradip Prajapati
//  FILE_NAME :- AHB_master_pkg.sv
//  EDITED_BY :- Pradip_Prajapati
//
//////////////////////////////////////////////////////////////////////////////////////////////////////////////

`include "ahb_master_agent_configuration.sv"
`include "ahb_master_transaction.sv"
`include "ahb_master_driver_callback.sv"
`include "ahb_master_driver_user_callback.sv"
`include "ahb_master_sequencer.sv"
`include "ahb_master_driver.sv"
`include "ahb_master_monitor.sv"
`include "ahb_master_checker.sv"
`include "ahb_master_agent.sv"
 
