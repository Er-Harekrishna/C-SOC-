//////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//  NAME      :- Pradip Prajapati
//  FILE_NAME :- AHB_slave_pkg.sv
//  EDITED_BY :- Pradip_Prajapati
//
//////////////////////////////////////////////////////////////////////////////////////////////////////////////

`include "ahb_slave_agent_configuration.sv"
`include "ahb_slave_transaction.sv"
`include "ahb_slave_driver_callback.sv"
`include "ahb_slave_driver_user_callback.sv"
`include "ahb_slave_sequencer.sv"
`include "ahb_slave_driver.sv"
`include "ahb_slave_monitor.sv"
//`include "AHB_slave_checker.sv"
`include "ahb_slave_agent.sv"

